module font_romtext(input[9:0] dx, dy,
							input win, lose,
							output on);
	
	logic [52:0] ROM1 [16];
	logic [61:0] ROM2 [16];
	logic [53:0] UP [16]; // W:UP
	logic [61:0] DOWN [16]; //S:DOWN
	logic [61:0] LEFT [16]; //A:LEFT
	logic [61:0] RIGHT [16]; //D:RIGHT
	logic [96:0] SetFlag [16]; //F:SET FLAG
	logic [102:0] ClearFlag [16]; //G:CLEAR FLAG
	logic [53:0] Clear [16]; //C:CLEAR
	
	
	always_comb
	begin
		if(dy < 17 & win & dx < 54) //win
			begin
				ROM1[0] = 53'b00000000000000000000000000000000000000000000000000000;
				ROM1[1] = 53'b00000000000000000000000000000000000000000000000000000;
				ROM1[2] = 53'b11000011001111100011000110001100001100011110011000110;
				ROM1[3] = 53'b11000011011000110011000110001100001100001100011100110;
				ROM1[4] = 53'b11000011011000110011000110001100001100001100011110110;
				ROM1[5] = 53'b11000011011000110011000110001100001100001100011111110;
				ROM1[6] = 53'b00111100011000110011000110001100001100001100011011110;
				ROM1[7] = 53'b00011000011000110011000110001101101100001100011001110;
				ROM1[8] = 53'b00011000011000110011000110001101101100001100011000110;
				ROM1[9] = 53'b00011000011000110011000110001111111100001100011000110;
			  ROM1[10] = 53'b00111000011000110011000110000110011000001100011000110;
			  ROM1[11] = 53'b00111100001111100001111100000110011000011110011000110;
			  ROM1[12] = 53'b00000000000000000000000000000000000000000000000000000;
			  ROM1[13] = 53'b00000000000000000000000000000000000000000000000000000;
			  ROM1[14] = 53'b00000000000000000000000000000000000000000000000000000;
			  ROM1[15] = 53'b00000000000000000000000000000000000000000000000000000;
				
				on = ROM1[dy][53-dx];
			end
		else if(dy < 17 & lose & dx < 64) //lose
		begin
			   ROM2[0] = 63'b000000000000000000000000000000000000000000000000000000000000000;
				ROM2[1] = 63'b000000000000000000000000000000000000000000000000000000000000000;
				ROM2[2] = 63'b110000110011111000110001100011110000001111100001111100011111110;
				ROM2[3] = 63'b110000110110001100110001100001100000011000110011000110001100110;
				ROM2[4] = 63'b110000110110001100110001100001100000011000110011000110001100010;
				ROM2[5] = 63'b110000110110001100110001100001100000011000110001100000001101000;
				ROM2[6] = 63'b001111000110001100110001100001100000011000110000111000001111000;
				ROM2[7] = 63'b000110000110001100110001100001100000011000110000001100001101000;
				ROM2[8] = 63'b000110000110001100110001100001100000011000110000000110001100000;
				ROM2[9] = 63'b000110000110001100110001100001100010011000110011000110001100010;
			  ROM2[10] = 63'b001110000110001100110001100001100110011000110011000110001100110;
			  ROM2[11] = 63'b001111000011111000011111000011111110001111100001111100011111110;
			  ROM2[12] = 63'b000000000000000000000000000000000000000000000000000000000000000;
			  ROM2[13] = 63'b000000000000000000000000000000000000000000000000000000000000000;
			  ROM2[14] = 63'b000000000000000000000000000000000000000000000000000000000000000;
			  ROM2[15] = 63'b000000000000000000000000000000000000000000000000000000000000000;
				
				on = ROM2[dy][63-dx];
		end
		else if(~win & ~lose & dy < 96 & dx < 35) // W:UP
		begin
			   UP[0] = 35'b00000000000000000000000000000000000;
				UP[1] = 35'b00000000000000000000000000000000000;
				UP[2] = 35'b00000000000000000011000110011111100;
				UP[3] = 35'b00000000000000000011000110001100110;
				UP[4] = 35'b11000011000011000011000110001100110;
				UP[5] = 35'b11000011000011000011000110001100110;
				UP[6] = 35'b11000011000000000011000110001111100;
				UP[7] = 35'b11011011000000000011000110001100000;
				UP[8] = 35'b11011011000000000011000110001100000;
				UP[9] = 35'b11111111000011000011000110001100000;
			  UP[10] = 35'b01100110000011000011000110001100000;
			  UP[11] = 35'b00000000000000000001111100011110000;
			  UP[12] = 35'b00000000000000000000000000000000000;
			  UP[13] = 35'b00000000000000000000000000000000000;
			  UP[14] = 35'b00000000000000000000000000000000000;
			  UP[15] = 35'b00000000000000000000000000000000000;
				
				on = UP[dy][35-dx];
		end
		else if(dy > 32 & dy > 96 & dy < 96+16 & dx < 53) //S:DOWN
		begin
			   DOWN[0] = 53'b0000000000000000000000000000000000000000000000000000;
				DOWN[1] = 53'b0000000000000000000000000000000000000000000000000000;
				DOWN[2] = 53'b1111100000000000111110000011111000110000110011000110;
				DOWN[3] = 53'b0110110000000000011011000110001100110000110011100110;
				DOWN[4] = 53'b0110011000011000011001100110001100110000110011110110;
				DOWN[5] = 53'b0110011000011000011001100110001100110000110011111110;
				DOWN[6] = 53'b0110011000000000011001100110001100110000110011011110;
				DOWN[7] = 53'b0110011000000000011001100110001100110110110011001110;
				DOWN[8] = 53'b0110011000000000011001100110001100110110110011000110;
				DOWN[9] = 53'b0110011000011000011001100110001100111111110011000110;
			  DOWN[10] = 53'b0110110000011000011011000110001100011001100011000110;
			  DOWN[11] = 53'b1111100000011000111110000011111000011001100011000110;
			  DOWN[12] = 53'b0000000000000000000000000000000000000000000000000000;
			  DOWN[13] = 53'b0000000000000000000000000000000000000000000000000000;
			  DOWN[14] = 53'b0000000000000000000000000000000000000000000000000000;
			  DOWN[15] = 53'b0000000000000000000000000000000000000000000000000000;
				
				on = DOWN[dy][53-dx];
		end
		else if(dy > 32 & dy > 96+16 & dy < 96+16+16 & dx < 54) //A:LEFT
		begin
			   LEFT[0] = 52'b0000000000000000000000000000000000000000000000000000;
				LEFT[1] = 52'b0000000000000000000000000000000000000000000000000000;
				LEFT[2] = 52'b0001000000000000011110000011111110011111110011111111;
				LEFT[3] = 52'b0011100000000000001100000001100110001100110011011011;
				LEFT[4] = 52'b0110110000001100001100000001100010001100010010011001;
				LEFT[5] = 52'b1100011000001100001100000001101000001101000000011000;
				LEFT[6] = 52'b1100011000000000001100000001111000001111000000011000;
				LEFT[7] = 52'b1111111000000000001100000001101000001101000000011000;
				LEFT[8] = 52'b1100011000000000001100000001100000001100000000011000;
				LEFT[9] = 52'b1100011000001100001100010001100010001100000000011000;
			  LEFT[10] = 52'b1100011000001100001100110001100110001100000000011000;
			  LEFT[11] = 52'b1100011000000000011111110011111110011110000000111100;
			  LEFT[12] = 52'b0000000000000000000000000000000000000000000000000000;
			  LEFT[13] = 52'b0000000000000000000000000000000000000000000000000000;
			  LEFT[14] = 52'b0000000000000000000000000000000000000000000000000000;
			  LEFT[15] = 52'b0000000000000000000000000000000000000000000000000000;
				
				on = LEFT[dy][54-dx];
		end
		else if(dy > 96+16+16 & dy < 96+16+16+16 & dx < 61) //D:RIGHT
		begin
			   RIGHT[0] = 61'b00000000000000000000000000000000000000000000000000000000000;
				RIGHT[1] = 61'b00000000000000000000000000000000000000000000000000000000000;
				RIGHT[2] = 61'b11111000000000001111110000011110000111100011000110011111111;
				RIGHT[3] = 61'b01101100000000000110011000001100001100110011000110011011011;
				RIGHT[4] = 61'b01100110000110000110011000001100011000010011000110010011001;
				RIGHT[5] = 61'b01100110000110000110011000001100011000000011000110000011000;
				RIGHT[6] = 61'b01100110000000000111110000001100011000000011111110000011000;
				RIGHT[7] = 61'b01100110000000000110110000001100011011110011000110000011000;
				RIGHT[8] = 61'b01100110000000000110011000001100011000110011000110000011000;
				RIGHT[9] = 61'b01100110000110000110011000001100011000110011000110000011000;
			  RIGHT[10] = 61'b01101100000110000110011000001100011000110011000110000011000;
			  RIGHT[11] = 61'b11111000000000001110011000011110001111100011000110000111100;
			  RIGHT[12] = 61'b00000000000000000000000000000000000000000000000000000000000;
			  RIGHT[13] = 61'b00000000000000000000000000000000000000000000000000000000000;
			  RIGHT[14] = 61'b00000000000000000000000000000000000000000000000000000000000;
			  RIGHT[15] = 61'b00000000000000000000000000000000000000000000000000000000000;
				
				on = RIGHT[dy][61-dx];
		end
		else if(dy > 96+16+16+16 & dy < 96+16+16+16+16 & dx < 96) //F:SET FLAG
		begin
			   SetFlag[0] = 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				SetFlag[1] = 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				SetFlag[2] = 96'b011111100000011000001111111000011111100011111111000000000111111000011000000000111000000111111000;
				SetFlag[3] = 96'b011000100000011000001100011000011000100010011001000000000110001000011000000001101100001100001000;
				SetFlag[4] = 96'b011000100000000000000110000000011010000000011000000000000110100000011000000011000110001100000000;
				SetFlag[5] = 96'b011010000000000000000011100000011110000000011000000000000111100000011000000011000110001100000000;
				SetFlag[6] = 96'b011110000000000000000000110000011010000000011000000000000110100000011000000011111110001101111000;
				SetFlag[7] = 96'b011010000000011000000000011000011000000000011000000000000110000000011000000011000110001100011000;
				SetFlag[8] = 96'b011000000000011000001100011000011000100000011000000000000110000000011000100011000110001100001100;
				SetFlag[9] = 96'b011000000000000000001100011000011001100000011000000000000110000000011001100011000110001100110000;
			  SetFlag[10] = 96'b111100000000000000000111110000111111100000111100000000001111000000111111100011000110000011110000;
			  SetFlag[11] = 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			  SetFlag[12] = 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			  SetFlag[13] = 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			  SetFlag[14] = 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			  SetFlag[15] = 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				
				on = SetFlag[dy][96-dx];
		end
		else if(dy > 96+16+16+16+16 & dy < 96+16+16+16+16+16 & dx < 102) //G:CLEAR FLAG
		begin
			   ClearFlag[0] = 102'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				ClearFlag[1] = 102'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				ClearFlag[2] = 102'b001111000000000000011110001111000011111110000010000111111000000000011111110011110000000010000000111100;
				ClearFlag[3] = 102'b011001100000000000110011000110000001100110000111000011001100000000001100110001100000000111000001100110;
				ClearFlag[4] = 102'b110000100000110001100001000110000001100010001101100011001100000000001100010001100000001101100011000010;
				ClearFlag[5] = 102'b110000000000110001100000000110000001101000011000110011001100000000001101000001100000011000110011000000;
				ClearFlag[6] = 102'b110000000000000001100000000110000001111000011000110011111000000000001111000001100000011000110011000000;
				ClearFlag[7] = 102'b110111100000000001100000000110000001101000011111110011011000000000001101000001100000011111110011011110;
				ClearFlag[8] = 102'b110001100000000001100000000110000001100000011000110011001100000000001100000001100000011000110011000110;
				ClearFlag[9] = 102'b110001100000110001100001000110001001100010011000110011001100000000001100000001100010011000110011000110;
			  ClearFlag[10] = 102'b011001100000110000110011000110011001100110011000110011001100000000001100000001100110011000110001100110;
			  ClearFlag[11] = 102'b001110100000000000011110001111111011111110011000110111001100000000011110000011111110011000110000111010;
			  ClearFlag[12] = 102'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			  ClearFlag[13] = 102'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			  ClearFlag[14] = 102'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			  ClearFlag[15] = 102'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				
				on = ClearFlag[dy][102-dx];
		end
		else if(dy > 96+16+16+16+16+16 & dy < 96+16+16+16+16+16+16 & dx < 53) //C:CLEAR
		begin
			   Clear[0] = 53'b0000000000000000000000000000000000000000000000000000;
				Clear[1] = 53'b0000000000000000000000000000000000000000000000000000;
				Clear[2] = 53'b0011110000000000001111000011111110000010000011111100;
				Clear[3] = 53'b0110011000000000011001100001100110000111000001100110;
				Clear[4] = 53'b1100001000001100110000100001100010001101100001100110;
				Clear[5] = 53'b1100000000001100110000000001101000011000110001100110;
				Clear[6] = 53'b1100000000000000110000000001111000011000110001111100;
				Clear[7] = 53'b1100000000000000110000000001101000011111110001101100;
				Clear[8] = 53'b1100000000000000110000000001100000011000110001100110;
				Clear[9] = 53'b1100001000001100110000100001100010011000110001100110;
			  Clear[10] = 53'b0110011000001100011001100001100110011000110001100110;
			  Clear[11] = 53'b0011110000000000001111000011111110011000110011100110;
			  Clear[12] = 53'b0000000000000000000000000000000000000000000000000000;
			  Clear[13] = 53'b0000000000000000000000000000000000000000000000000000;
			  Clear[14] = 53'b0000000000000000000000000000000000000000000000000000;
			  Clear[15] = 53'b0000000000000000000000000000000000000000000000000000;
				
				on = Clear[dy][53-dx];
		end
		else
			on = 1'b0;
	end
endmodule
