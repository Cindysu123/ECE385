module reg_3
(	
					input logic Clk, Reset, Load,
					input logic [2:0] D,
					output logic [2:0] Data_Out
);

always_ff @(posedge Clk or posedge Reset)
	begin
		if (Reset)
			Data_Out <= 3'b000;
		else if (Load)
			Data_Out <= D;
//		else if (Shift_En)
//		begin
//			Data_Out <= { Shift_In, Data_Out[2:1] };
//		end
	end
		
//		assign Shift_Out = Data_Out[0];
		
		
endmodule
